`timescale 1ns/1ps

module decoder_a(

    input a, b, c,
    output z0, z1, z2, z3, z4, z5, z6, z7

);

    assign z0 = (~a & ~b & ~c);
    assign z1 = (a & ~b & ~c);
    assign z2 = (~a & b & ~c);
    assign z3 = (a & b & ~c);
    assign z4 = (~a & ~b & c);
    assign z5 = (a & ~b & c);
    assign z6 = (~a & b & c);
    assign z7 = (a & b & c);

endmodule